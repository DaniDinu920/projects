`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   12:00:09 12/12/2020
// Design Name:   rail_fence
// Module Name:   C:/verilog/rail_fence/rail_test.v
// Project Name:  rail_fence
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: rail_fence
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module rail_test;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	rail_fence uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

